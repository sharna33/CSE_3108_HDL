// 2003009

module subOne(
  input wire [4:0] i,
  output wire [4:0] o
);
  assign o = i - 1;
endmodule