`timescale 1ns/1ps

module enc_case_tb;
    reg [3:0] Y;
    wire [3:0] A;

    enc_case uut(
        .Y(Y),
        .A(A)
    );

    initial begin
        $dumpfile("enc_case_tb.vcd");
        $dumpvars(0, enc_case_tb);
        
        Y[3] = 0; Y[2] = 0; Y[1] = 0; Y[0] = 0;
        #20;
    
        Y[3] = 0; Y[2] = 0; Y[1] = 0; Y[0] = 1;
        #20;

        Y[3] = 0; Y[2] = 0; Y[1] = 1; Y[0] = 0;
        #20;

        Y[3] = 0; Y[2] = 0; Y[1] = 1; Y[0] = 1;
        #20;

        Y[3] = 0; Y[2] = 1; Y[1] = 0; Y[0] = 0;
        #20;

        Y[3] = 0; Y[2] = 1; Y[1] = 0; Y[0] = 1;
        #20;

        Y[3] = 0; Y[2] = 1; Y[1] = 1; Y[0] = 0;
        #20;

        Y[3] = 0; Y[2] = 1; Y[1] = 1; Y[0] = 1;
        #20;

        Y[3] = 1; Y[2] = 0; Y[1] = 0; Y[0] = 0;
        #20;

        Y[3] = 1; Y[2] = 0; Y[1] = 0; Y[0] = 1;
        #20;

        Y[3] = 1; Y[2] = 0; Y[1] = 1; Y[0] = 0;
        #20;

        Y[3] = 1; Y[2] = 0; Y[1] = 1; Y[0] = 1;
        #20;

        Y[3] = 1; Y[2] = 1; Y[1] = 0; Y[0] = 0;
        #20;

        Y[3] = 1; Y[2] = 1; Y[1] = 0; Y[0] = 1; 
        #20;

        Y[3] = 1; Y[2] = 1; Y[1] = 1; Y[0] = 0;
        #20;

        Y[3] = 1; Y[2] = 1; Y[1] = 1; Y[0] = 1;
        #20;

        $finish;
    end

    initial begin
        $monitor("Y = %b, A = %b", Y, A);
    end

endmodule